module FourToOneMux(LEDR, SW);
	input [9:0] SW;
	output [9:8] LEDR;
	
	
endmodule 